magic
tech sky130A
timestamp 1716270487
<< nwell >>
rect -100 -150 450 300
<< nmos >>
rect 45 -450 60 -350
rect 295 -450 310 -350
<< pmos >>
rect 45 -100 60 100
rect 295 -100 310 100
<< ndiff >>
rect 5 -365 45 -350
rect 5 -430 10 -365
rect 35 -430 45 -365
rect 5 -450 45 -430
rect 60 -365 100 -350
rect 60 -430 70 -365
rect 95 -430 100 -365
rect 60 -450 100 -430
rect 255 -365 295 -350
rect 255 -430 260 -365
rect 285 -430 295 -365
rect 255 -450 295 -430
rect 310 -365 350 -350
rect 310 -430 320 -365
rect 345 -430 350 -365
rect 310 -450 350 -430
<< pdiff >>
rect -40 85 45 100
rect -40 -90 -30 85
rect 30 -90 45 85
rect -40 -100 45 -90
rect 60 85 145 100
rect 60 -90 75 85
rect 135 -90 145 85
rect 60 -100 145 -90
rect 210 85 295 100
rect 210 -90 220 85
rect 280 -90 295 85
rect 210 -100 295 -90
rect 310 85 395 100
rect 310 -90 325 85
rect 385 -90 395 85
rect 310 -100 395 -90
<< ndiffc >>
rect 10 -430 35 -365
rect 70 -430 95 -365
rect 260 -430 285 -365
rect 320 -430 345 -365
<< pdiffc >>
rect -30 -90 30 85
rect 75 -90 135 85
rect 220 -90 280 85
rect 325 -90 385 85
<< psubdiff >>
rect 85 -535 230 -520
rect 85 -560 105 -535
rect 215 -560 230 -535
rect 85 -575 230 -560
<< nsubdiff >>
rect 50 235 300 250
rect 50 170 85 235
rect 275 170 300 235
rect 50 150 300 170
<< psubdiffcont >>
rect 105 -560 215 -535
<< nsubdiffcont >>
rect 85 170 275 235
<< poly >>
rect 45 100 60 115
rect 295 100 310 115
rect 45 -240 60 -100
rect -25 -250 60 -240
rect -25 -270 -15 -250
rect 25 -270 60 -250
rect -25 -285 60 -270
rect 45 -350 60 -285
rect 295 -240 310 -100
rect 295 -250 380 -240
rect 295 -270 325 -250
rect 365 -270 380 -250
rect 295 -285 380 -270
rect 295 -350 310 -285
rect 45 -500 60 -450
rect 295 -500 310 -450
<< polycont >>
rect -15 -270 25 -250
rect 325 -270 365 -250
<< locali >>
rect 50 235 300 250
rect 50 175 85 235
rect -20 170 85 175
rect 275 170 300 235
rect -20 150 300 170
rect -20 100 0 150
rect 220 100 240 150
rect -40 85 40 100
rect -40 -90 -30 85
rect 30 -90 40 85
rect -40 -100 40 -90
rect 65 85 145 100
rect 65 -90 75 85
rect 135 -90 145 85
rect 65 -100 145 -90
rect 210 85 290 100
rect 210 -90 220 85
rect 280 -90 290 85
rect 210 -100 290 -90
rect 315 85 395 100
rect 315 -90 325 85
rect 385 -90 395 85
rect 315 -100 395 -90
rect 80 -151 125 -100
rect 326 -149 368 -100
rect 201 -151 368 -149
rect 80 -163 368 -151
rect 80 -200 370 -163
rect -25 -250 45 -240
rect -25 -270 -15 -250
rect 25 -270 45 -250
rect -25 -285 45 -270
rect 80 -350 100 -200
rect 310 -250 380 -240
rect 310 -270 325 -250
rect 365 -270 380 -250
rect 310 -285 380 -270
rect 5 -365 40 -350
rect 5 -430 10 -365
rect 35 -430 40 -365
rect 5 -450 40 -430
rect 65 -365 100 -350
rect 65 -430 70 -365
rect 95 -430 100 -365
rect 65 -450 100 -430
rect 255 -365 290 -350
rect 255 -430 260 -365
rect 285 -430 290 -365
rect 255 -450 290 -430
rect 315 -365 350 -350
rect 315 -430 320 -365
rect 345 -430 350 -365
rect 315 -450 350 -430
rect 255 -520 275 -450
rect 85 -535 275 -520
rect 85 -560 105 -535
rect 215 -540 275 -535
rect 215 -560 230 -540
rect 85 -575 230 -560
<< viali >>
rect 85 170 275 235
rect -15 -270 25 -250
rect 325 -270 365 -250
rect 10 -430 35 -365
rect 320 -430 345 -365
rect 105 -560 215 -535
<< metal1 >>
rect 50 235 300 250
rect 50 170 85 235
rect 275 170 300 235
rect 50 150 300 170
rect -25 -250 45 -240
rect -25 -270 -15 -250
rect 25 -270 45 -250
rect -25 -285 45 -270
rect 310 -250 380 -240
rect 310 -270 325 -250
rect 365 -270 380 -250
rect 310 -285 380 -270
rect 5 -365 350 -350
rect 5 -430 10 -365
rect 35 -375 320 -365
rect 35 -430 40 -375
rect 5 -450 40 -430
rect 315 -430 320 -375
rect 345 -430 350 -365
rect 315 -450 350 -430
rect 85 -535 230 -520
rect 85 -560 105 -535
rect 215 -560 230 -535
rect 85 -575 230 -560
<< labels >>
rlabel metal1 -20 -260 -20 -260 1 A
port 1 n
rlabel metal1 370 -260 370 -260 1 B
port 2 n
rlabel metal1 200 -530 200 -530 1 gnd
port 3 n
rlabel metal1 245 240 245 240 1 vdd
port 4 n
<< end >>
