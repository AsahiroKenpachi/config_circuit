magic
tech sky130A
timestamp 1716356529
<< nwell >>
rect -100 -150 1715 300
rect -100 -1100 1705 -650
rect -100 -2095 1105 -1645
rect 1255 -2095 1765 -1645
<< nmos >>
rect 45 -450 60 -350
rect 295 -450 310 -350
rect 795 -450 810 -350
rect 1045 -450 1060 -350
rect 1310 -450 1325 -350
rect 45 -1400 60 -1300
rect 295 -1400 310 -1300
rect 780 -1400 795 -1300
rect 1030 -1400 1045 -1300
rect 1300 -1400 1315 -1300
rect 30 -2395 45 -2295
rect 280 -2395 295 -2295
rect 700 -2395 715 -2295
rect 950 -2395 965 -2295
rect 1360 -2395 1375 -2295
<< pmos >>
rect 45 -100 60 100
rect 295 -100 310 100
rect 795 -100 810 100
rect 1045 -100 1060 100
rect 1310 -100 1325 100
rect 45 -1050 60 -850
rect 295 -1050 310 -850
rect 780 -1050 795 -850
rect 1030 -1050 1045 -850
rect 1300 -1050 1315 -850
rect 30 -2045 45 -1845
rect 280 -2045 295 -1845
rect 700 -2045 715 -1845
rect 950 -2045 965 -1845
rect 1360 -2045 1375 -1845
<< ndiff >>
rect 5 -365 45 -350
rect 5 -430 10 -365
rect 35 -430 45 -365
rect 5 -450 45 -430
rect 60 -365 100 -350
rect 60 -430 70 -365
rect 95 -430 100 -365
rect 60 -450 100 -430
rect 255 -365 295 -350
rect 255 -430 260 -365
rect 285 -430 295 -365
rect 255 -450 295 -430
rect 310 -365 350 -350
rect 310 -430 320 -365
rect 345 -430 350 -365
rect 310 -450 350 -430
rect 755 -365 795 -350
rect 755 -430 760 -365
rect 785 -430 795 -365
rect 755 -450 795 -430
rect 810 -365 850 -350
rect 810 -430 820 -365
rect 845 -430 850 -365
rect 810 -450 850 -430
rect 1005 -365 1045 -350
rect 1005 -430 1010 -365
rect 1035 -430 1045 -365
rect 1005 -450 1045 -430
rect 1060 -365 1100 -350
rect 1060 -430 1070 -365
rect 1095 -430 1100 -365
rect 1060 -450 1100 -430
rect 1270 -365 1310 -350
rect 1270 -430 1275 -365
rect 1300 -430 1310 -365
rect 1270 -450 1310 -430
rect 1325 -365 1365 -350
rect 1325 -430 1335 -365
rect 1360 -430 1365 -365
rect 1325 -450 1365 -430
rect 5 -1315 45 -1300
rect 5 -1380 10 -1315
rect 35 -1380 45 -1315
rect 5 -1400 45 -1380
rect 60 -1315 100 -1300
rect 60 -1380 70 -1315
rect 95 -1380 100 -1315
rect 60 -1400 100 -1380
rect 255 -1315 295 -1300
rect 255 -1380 260 -1315
rect 285 -1380 295 -1315
rect 255 -1400 295 -1380
rect 310 -1315 350 -1300
rect 310 -1380 320 -1315
rect 345 -1380 350 -1315
rect 310 -1400 350 -1380
rect 740 -1315 780 -1300
rect 740 -1380 745 -1315
rect 770 -1380 780 -1315
rect 740 -1400 780 -1380
rect 795 -1315 835 -1300
rect 795 -1380 805 -1315
rect 830 -1380 835 -1315
rect 795 -1400 835 -1380
rect 990 -1315 1030 -1300
rect 990 -1380 995 -1315
rect 1020 -1380 1030 -1315
rect 990 -1400 1030 -1380
rect 1045 -1315 1085 -1300
rect 1045 -1380 1055 -1315
rect 1080 -1380 1085 -1315
rect 1045 -1400 1085 -1380
rect 1260 -1315 1300 -1300
rect 1260 -1380 1265 -1315
rect 1290 -1380 1300 -1315
rect 1260 -1400 1300 -1380
rect 1315 -1315 1355 -1300
rect 1315 -1380 1325 -1315
rect 1350 -1380 1355 -1315
rect 1315 -1400 1355 -1380
rect -10 -2310 30 -2295
rect -10 -2375 -5 -2310
rect 20 -2375 30 -2310
rect -10 -2395 30 -2375
rect 45 -2310 85 -2295
rect 45 -2375 55 -2310
rect 80 -2375 85 -2310
rect 45 -2395 85 -2375
rect 240 -2310 280 -2295
rect 240 -2375 245 -2310
rect 270 -2375 280 -2310
rect 240 -2395 280 -2375
rect 295 -2310 335 -2295
rect 295 -2375 305 -2310
rect 330 -2375 335 -2310
rect 295 -2395 335 -2375
rect 660 -2310 700 -2295
rect 660 -2375 665 -2310
rect 690 -2375 700 -2310
rect 660 -2395 700 -2375
rect 715 -2310 755 -2295
rect 715 -2375 725 -2310
rect 750 -2375 755 -2310
rect 715 -2395 755 -2375
rect 910 -2310 950 -2295
rect 910 -2375 915 -2310
rect 940 -2375 950 -2310
rect 910 -2395 950 -2375
rect 965 -2310 1005 -2295
rect 965 -2375 975 -2310
rect 1000 -2375 1005 -2310
rect 965 -2395 1005 -2375
rect 1320 -2310 1360 -2295
rect 1320 -2375 1325 -2310
rect 1350 -2375 1360 -2310
rect 1320 -2395 1360 -2375
rect 1375 -2310 1415 -2295
rect 1375 -2375 1385 -2310
rect 1410 -2375 1415 -2310
rect 1375 -2395 1415 -2375
<< pdiff >>
rect -40 85 45 100
rect -40 -90 -30 85
rect 30 -90 45 85
rect -40 -100 45 -90
rect 60 85 145 100
rect 60 -90 75 85
rect 135 -90 145 85
rect 60 -100 145 -90
rect 210 85 295 100
rect 210 -90 220 85
rect 280 -90 295 85
rect 210 -100 295 -90
rect 310 85 395 100
rect 310 -90 325 85
rect 385 -90 395 85
rect 310 -100 395 -90
rect 710 85 795 100
rect 710 -90 720 85
rect 780 -90 795 85
rect 710 -100 795 -90
rect 810 85 895 100
rect 810 -90 825 85
rect 885 -90 895 85
rect 810 -100 895 -90
rect 960 85 1045 100
rect 960 -90 970 85
rect 1030 -90 1045 85
rect 960 -100 1045 -90
rect 1060 85 1145 100
rect 1060 -90 1075 85
rect 1135 -90 1145 85
rect 1060 -100 1145 -90
rect 1225 85 1310 100
rect 1225 -90 1235 85
rect 1295 -90 1310 85
rect 1225 -100 1310 -90
rect 1325 85 1410 100
rect 1325 -90 1340 85
rect 1400 -90 1410 85
rect 1325 -100 1410 -90
rect -40 -865 45 -850
rect -40 -1040 -30 -865
rect 30 -1040 45 -865
rect -40 -1050 45 -1040
rect 60 -865 145 -850
rect 60 -1040 75 -865
rect 135 -1040 145 -865
rect 60 -1050 145 -1040
rect 210 -865 295 -850
rect 210 -1040 220 -865
rect 280 -1040 295 -865
rect 210 -1050 295 -1040
rect 310 -865 395 -850
rect 310 -1040 325 -865
rect 385 -1040 395 -865
rect 310 -1050 395 -1040
rect 695 -865 780 -850
rect 695 -1040 705 -865
rect 765 -1040 780 -865
rect 695 -1050 780 -1040
rect 795 -865 880 -850
rect 795 -1040 810 -865
rect 870 -1040 880 -865
rect 795 -1050 880 -1040
rect 945 -865 1030 -850
rect 945 -1040 955 -865
rect 1015 -1040 1030 -865
rect 945 -1050 1030 -1040
rect 1045 -865 1130 -850
rect 1045 -1040 1060 -865
rect 1120 -1040 1130 -865
rect 1045 -1050 1130 -1040
rect 1215 -865 1300 -850
rect 1215 -1040 1225 -865
rect 1285 -1040 1300 -865
rect 1215 -1050 1300 -1040
rect 1315 -865 1400 -850
rect 1315 -1040 1330 -865
rect 1390 -1040 1400 -865
rect 1315 -1050 1400 -1040
rect -55 -1860 30 -1845
rect -55 -2035 -45 -1860
rect 15 -2035 30 -1860
rect -55 -2045 30 -2035
rect 45 -1860 130 -1845
rect 45 -2035 60 -1860
rect 120 -2035 130 -1860
rect 45 -2045 130 -2035
rect 195 -1860 280 -1845
rect 195 -2035 205 -1860
rect 265 -2035 280 -1860
rect 195 -2045 280 -2035
rect 295 -1860 380 -1845
rect 295 -2035 310 -1860
rect 370 -2035 380 -1860
rect 295 -2045 380 -2035
rect 615 -1860 700 -1845
rect 615 -2035 625 -1860
rect 685 -2035 700 -1860
rect 615 -2045 700 -2035
rect 715 -1860 800 -1845
rect 715 -2035 730 -1860
rect 790 -2035 800 -1860
rect 715 -2045 800 -2035
rect 865 -1860 950 -1845
rect 865 -2035 875 -1860
rect 935 -2035 950 -1860
rect 865 -2045 950 -2035
rect 965 -1860 1050 -1845
rect 965 -2035 980 -1860
rect 1040 -2035 1050 -1860
rect 965 -2045 1050 -2035
rect 1275 -1860 1360 -1845
rect 1275 -2035 1285 -1860
rect 1345 -2035 1360 -1860
rect 1275 -2045 1360 -2035
rect 1375 -1860 1460 -1845
rect 1375 -2035 1390 -1860
rect 1450 -2035 1460 -1860
rect 1375 -2045 1460 -2035
<< ndiffc >>
rect 10 -430 35 -365
rect 70 -430 95 -365
rect 260 -430 285 -365
rect 320 -430 345 -365
rect 760 -430 785 -365
rect 820 -430 845 -365
rect 1010 -430 1035 -365
rect 1070 -430 1095 -365
rect 1275 -430 1300 -365
rect 1335 -430 1360 -365
rect 10 -1380 35 -1315
rect 70 -1380 95 -1315
rect 260 -1380 285 -1315
rect 320 -1380 345 -1315
rect 745 -1380 770 -1315
rect 805 -1380 830 -1315
rect 995 -1380 1020 -1315
rect 1055 -1380 1080 -1315
rect 1265 -1380 1290 -1315
rect 1325 -1380 1350 -1315
rect -5 -2375 20 -2310
rect 55 -2375 80 -2310
rect 245 -2375 270 -2310
rect 305 -2375 330 -2310
rect 665 -2375 690 -2310
rect 725 -2375 750 -2310
rect 915 -2375 940 -2310
rect 975 -2375 1000 -2310
rect 1325 -2375 1350 -2310
rect 1385 -2375 1410 -2310
<< pdiffc >>
rect -30 -90 30 85
rect 75 -90 135 85
rect 220 -90 280 85
rect 325 -90 385 85
rect 720 -90 780 85
rect 825 -90 885 85
rect 970 -90 1030 85
rect 1075 -90 1135 85
rect 1235 -90 1295 85
rect 1340 -90 1400 85
rect -30 -1040 30 -865
rect 75 -1040 135 -865
rect 220 -1040 280 -865
rect 325 -1040 385 -865
rect 705 -1040 765 -865
rect 810 -1040 870 -865
rect 955 -1040 1015 -865
rect 1060 -1040 1120 -865
rect 1225 -1040 1285 -865
rect 1330 -1040 1390 -865
rect -45 -2035 15 -1860
rect 60 -2035 120 -1860
rect 205 -2035 265 -1860
rect 310 -2035 370 -1860
rect 625 -2035 685 -1860
rect 730 -2035 790 -1860
rect 875 -2035 935 -1860
rect 980 -2035 1040 -1860
rect 1285 -2035 1345 -1860
rect 1390 -2035 1450 -1860
<< psubdiff >>
rect 85 -535 230 -520
rect 85 -560 105 -535
rect 215 -560 230 -535
rect 85 -575 230 -560
rect 835 -535 980 -520
rect 835 -560 855 -535
rect 965 -560 980 -535
rect 835 -575 980 -560
rect 1350 -535 1495 -520
rect 1350 -560 1370 -535
rect 1480 -560 1495 -535
rect 1350 -575 1495 -560
rect 85 -1485 230 -1470
rect 85 -1510 105 -1485
rect 215 -1510 230 -1485
rect 85 -1525 230 -1510
rect 820 -1485 965 -1470
rect 820 -1510 840 -1485
rect 950 -1510 965 -1485
rect 820 -1525 965 -1510
rect 1340 -1485 1485 -1470
rect 1340 -1510 1360 -1485
rect 1470 -1510 1485 -1485
rect 1340 -1525 1485 -1510
rect 70 -2480 215 -2465
rect 70 -2505 90 -2480
rect 200 -2505 215 -2480
rect 70 -2520 215 -2505
rect 740 -2480 885 -2465
rect 740 -2505 760 -2480
rect 870 -2505 885 -2480
rect 740 -2520 885 -2505
rect 1400 -2480 1545 -2465
rect 1400 -2505 1420 -2480
rect 1530 -2505 1545 -2480
rect 1400 -2520 1545 -2505
<< nsubdiff >>
rect 50 235 300 250
rect 50 170 85 235
rect 275 170 300 235
rect 50 150 300 170
rect 800 235 1050 250
rect 800 170 835 235
rect 1025 170 1050 235
rect 800 150 1050 170
rect 1315 235 1565 250
rect 1315 170 1350 235
rect 1540 170 1565 235
rect 1315 150 1565 170
rect 50 -715 300 -700
rect 50 -780 85 -715
rect 275 -780 300 -715
rect 50 -800 300 -780
rect 785 -715 1035 -700
rect 785 -780 820 -715
rect 1010 -780 1035 -715
rect 785 -800 1035 -780
rect 1305 -715 1555 -700
rect 1305 -780 1340 -715
rect 1530 -780 1555 -715
rect 1305 -800 1555 -780
rect 35 -1710 285 -1695
rect 35 -1775 70 -1710
rect 260 -1775 285 -1710
rect 35 -1795 285 -1775
rect 705 -1710 955 -1695
rect 705 -1775 740 -1710
rect 930 -1775 955 -1710
rect 705 -1795 955 -1775
rect 1365 -1710 1615 -1695
rect 1365 -1775 1400 -1710
rect 1590 -1775 1615 -1710
rect 1365 -1795 1615 -1775
<< psubdiffcont >>
rect 105 -560 215 -535
rect 855 -560 965 -535
rect 1370 -560 1480 -535
rect 105 -1510 215 -1485
rect 840 -1510 950 -1485
rect 1360 -1510 1470 -1485
rect 90 -2505 200 -2480
rect 760 -2505 870 -2480
rect 1420 -2505 1530 -2480
<< nsubdiffcont >>
rect 85 170 275 235
rect 835 170 1025 235
rect 1350 170 1540 235
rect 85 -780 275 -715
rect 820 -780 1010 -715
rect 1340 -780 1530 -715
rect 70 -1775 260 -1710
rect 740 -1775 930 -1710
rect 1400 -1775 1590 -1710
<< poly >>
rect 45 100 60 115
rect 295 100 310 115
rect 795 100 810 115
rect 1045 100 1060 115
rect 1310 100 1325 115
rect 45 -240 60 -100
rect -25 -250 60 -240
rect -25 -270 -15 -250
rect 25 -270 60 -250
rect -25 -285 60 -270
rect 45 -350 60 -285
rect 295 -240 310 -100
rect 365 -160 440 -145
rect 365 -180 380 -160
rect 425 -180 440 -160
rect 365 -200 440 -180
rect 795 -240 810 -100
rect 295 -250 380 -240
rect 295 -270 325 -250
rect 365 -270 380 -250
rect 295 -285 380 -270
rect 725 -250 810 -240
rect 725 -270 735 -250
rect 775 -270 810 -250
rect 725 -285 810 -270
rect 295 -350 310 -285
rect 795 -350 810 -285
rect 1045 -240 1060 -100
rect 1095 -150 1165 -135
rect 1095 -170 1110 -150
rect 1155 -170 1165 -150
rect 1095 -190 1165 -170
rect 1310 -240 1325 -100
rect 1365 -175 1435 -160
rect 1365 -195 1380 -175
rect 1420 -195 1435 -175
rect 1365 -215 1435 -195
rect 1045 -250 1130 -240
rect 1045 -270 1075 -250
rect 1115 -270 1130 -250
rect 1045 -285 1130 -270
rect 1240 -250 1325 -240
rect 1240 -270 1250 -250
rect 1290 -270 1325 -250
rect 1240 -285 1325 -270
rect 1045 -350 1060 -285
rect 1310 -350 1325 -285
rect 45 -500 60 -450
rect 295 -500 310 -450
rect 795 -500 810 -450
rect 1045 -500 1060 -450
rect 1310 -500 1325 -450
rect 45 -850 60 -835
rect 295 -850 310 -835
rect 780 -850 795 -835
rect 1030 -850 1045 -835
rect 1300 -850 1315 -835
rect 45 -1190 60 -1050
rect -25 -1200 60 -1190
rect -25 -1220 -15 -1200
rect 25 -1220 60 -1200
rect -25 -1235 60 -1220
rect 45 -1300 60 -1235
rect 295 -1190 310 -1050
rect 365 -1110 435 -1095
rect 365 -1130 380 -1110
rect 420 -1130 435 -1110
rect 365 -1150 435 -1130
rect 780 -1190 795 -1050
rect 295 -1200 380 -1190
rect 295 -1220 325 -1200
rect 365 -1220 380 -1200
rect 295 -1235 380 -1220
rect 710 -1200 795 -1190
rect 710 -1220 720 -1200
rect 760 -1220 795 -1200
rect 710 -1235 795 -1220
rect 295 -1300 310 -1235
rect 780 -1300 795 -1235
rect 1030 -1190 1045 -1050
rect 1075 -1115 1145 -1100
rect 1075 -1135 1090 -1115
rect 1130 -1135 1145 -1115
rect 1075 -1155 1145 -1135
rect 1300 -1190 1315 -1050
rect 1355 -1115 1425 -1100
rect 1355 -1135 1370 -1115
rect 1410 -1135 1425 -1115
rect 1355 -1155 1425 -1135
rect 1030 -1200 1115 -1190
rect 1030 -1220 1060 -1200
rect 1100 -1220 1115 -1200
rect 1030 -1235 1115 -1220
rect 1230 -1200 1315 -1190
rect 1230 -1220 1240 -1200
rect 1280 -1220 1315 -1200
rect 1230 -1235 1315 -1220
rect 1030 -1300 1045 -1235
rect 1300 -1300 1315 -1235
rect 45 -1450 60 -1400
rect 295 -1450 310 -1400
rect 780 -1450 795 -1400
rect 1030 -1450 1045 -1400
rect 1300 -1450 1315 -1400
rect 30 -1845 45 -1830
rect 280 -1845 295 -1830
rect 700 -1845 715 -1830
rect 950 -1845 965 -1830
rect 1360 -1845 1375 -1830
rect 30 -2185 45 -2045
rect -40 -2195 45 -2185
rect -40 -2215 -30 -2195
rect 10 -2215 45 -2195
rect -40 -2230 45 -2215
rect 30 -2295 45 -2230
rect 280 -2185 295 -2045
rect 325 -2110 395 -2095
rect 325 -2130 340 -2110
rect 380 -2130 395 -2110
rect 325 -2150 395 -2130
rect 700 -2185 715 -2045
rect 280 -2195 365 -2185
rect 280 -2215 310 -2195
rect 350 -2215 365 -2195
rect 280 -2230 365 -2215
rect 630 -2195 715 -2185
rect 630 -2215 640 -2195
rect 680 -2215 715 -2195
rect 630 -2230 715 -2215
rect 280 -2295 295 -2230
rect 700 -2295 715 -2230
rect 950 -2185 965 -2045
rect 1020 -2105 1090 -2100
rect 1020 -2125 1035 -2105
rect 1075 -2125 1090 -2105
rect 1020 -2145 1090 -2125
rect 1360 -2185 1375 -2045
rect 1415 -2125 1485 -2110
rect 1415 -2145 1430 -2125
rect 1470 -2145 1485 -2125
rect 1415 -2165 1485 -2145
rect 950 -2195 1035 -2185
rect 950 -2215 980 -2195
rect 1020 -2215 1035 -2195
rect 950 -2230 1035 -2215
rect 1290 -2195 1375 -2185
rect 1290 -2215 1300 -2195
rect 1340 -2215 1375 -2195
rect 1290 -2230 1375 -2215
rect 950 -2295 965 -2230
rect 1360 -2295 1375 -2230
rect 30 -2445 45 -2395
rect 280 -2445 295 -2395
rect 700 -2445 715 -2395
rect 950 -2445 965 -2395
rect 1360 -2445 1375 -2395
<< polycont >>
rect -15 -270 25 -250
rect 380 -180 425 -160
rect 325 -270 365 -250
rect 735 -270 775 -250
rect 1110 -170 1155 -150
rect 1380 -195 1420 -175
rect 1075 -270 1115 -250
rect 1250 -270 1290 -250
rect -15 -1220 25 -1200
rect 380 -1130 420 -1110
rect 325 -1220 365 -1200
rect 720 -1220 760 -1200
rect 1090 -1135 1130 -1115
rect 1370 -1135 1410 -1115
rect 1060 -1220 1100 -1200
rect 1240 -1220 1280 -1200
rect -30 -2215 10 -2195
rect 340 -2130 380 -2110
rect 310 -2215 350 -2195
rect 640 -2215 680 -2195
rect 1035 -2125 1075 -2105
rect 1430 -2145 1470 -2125
rect 980 -2215 1020 -2195
rect 1300 -2215 1340 -2195
<< locali >>
rect 50 235 300 250
rect 50 175 85 235
rect -20 170 85 175
rect 275 170 300 235
rect 800 235 1050 250
rect 800 175 835 235
rect -20 150 300 170
rect 730 170 835 175
rect 1025 170 1050 235
rect 1315 235 1565 250
rect 1315 175 1350 235
rect 730 150 1050 170
rect 1245 170 1350 175
rect 1540 170 1565 235
rect 1245 150 1565 170
rect -20 100 0 150
rect 220 100 240 150
rect 730 100 750 150
rect 1245 100 1265 150
rect -40 85 40 100
rect -40 -90 -30 85
rect 30 -90 40 85
rect -40 -100 40 -90
rect 65 85 145 100
rect 65 -90 75 85
rect 135 -90 145 85
rect 65 -100 145 -90
rect 210 85 290 100
rect 210 -90 220 85
rect 280 -90 290 85
rect 210 -100 290 -90
rect 315 85 395 100
rect 315 -90 325 85
rect 385 -90 395 85
rect 315 -100 395 -90
rect 710 85 790 100
rect 710 -90 720 85
rect 780 -90 790 85
rect 710 -100 790 -90
rect 815 95 895 100
rect 960 95 1040 100
rect 815 85 1040 95
rect 815 -90 825 85
rect 885 45 970 85
rect 885 -90 895 45
rect 815 -100 895 -90
rect 960 -90 970 45
rect 1030 -90 1040 85
rect 960 -100 1040 -90
rect 1065 85 1145 100
rect 1065 -90 1075 85
rect 1135 -90 1145 85
rect 1065 -100 1145 -90
rect 1225 85 1305 100
rect 1225 -90 1235 85
rect 1295 -90 1305 85
rect 1225 -100 1305 -90
rect 1330 85 1410 100
rect 1330 -90 1340 85
rect 1400 -90 1410 85
rect 1330 -100 1410 -90
rect 80 -151 125 -100
rect 326 -145 368 -100
rect 1090 -120 1130 -100
rect 885 -135 1130 -120
rect 326 -149 610 -145
rect 201 -151 610 -149
rect 80 -160 610 -151
rect 80 -180 380 -160
rect 425 -180 610 -160
rect 80 -200 610 -180
rect -25 -250 45 -240
rect -25 -270 -15 -250
rect 25 -270 45 -250
rect -25 -285 45 -270
rect 80 -350 100 -200
rect 310 -250 435 -240
rect 310 -270 325 -250
rect 365 -270 435 -250
rect 310 -285 435 -270
rect 5 -365 40 -350
rect 5 -430 10 -365
rect 35 -430 40 -365
rect 5 -450 40 -430
rect 65 -365 100 -350
rect 65 -430 70 -365
rect 95 -430 100 -365
rect 65 -450 100 -430
rect 255 -365 290 -350
rect 255 -430 260 -365
rect 285 -430 290 -365
rect 255 -450 290 -430
rect 315 -365 350 -350
rect 315 -430 320 -365
rect 345 -430 350 -365
rect 315 -450 350 -430
rect 255 -520 275 -450
rect 85 -535 275 -520
rect 85 -560 105 -535
rect 215 -540 275 -535
rect 215 -560 230 -540
rect 85 -575 230 -560
rect 405 -595 435 -285
rect -175 -630 435 -595
rect -175 -1190 -105 -630
rect 50 -715 300 -700
rect 50 -775 85 -715
rect -20 -780 85 -775
rect 275 -780 300 -715
rect -20 -800 300 -780
rect -20 -850 0 -800
rect 220 -850 240 -800
rect -40 -865 40 -850
rect -40 -1040 -30 -865
rect 30 -1040 40 -865
rect -40 -1050 40 -1040
rect 65 -865 145 -850
rect 65 -1040 75 -865
rect 135 -1040 145 -865
rect 65 -1050 145 -1040
rect 210 -865 290 -850
rect 210 -1040 220 -865
rect 280 -1040 290 -865
rect 210 -1050 290 -1040
rect 315 -865 395 -850
rect 315 -1040 325 -865
rect 385 -1040 395 -865
rect 315 -1050 395 -1040
rect 80 -1101 125 -1050
rect 326 -1095 368 -1050
rect 326 -1099 450 -1095
rect 201 -1101 450 -1099
rect 80 -1110 450 -1101
rect 80 -1130 380 -1110
rect 420 -1130 450 -1110
rect 80 -1150 450 -1130
rect -175 -1200 45 -1190
rect -175 -1220 -15 -1200
rect 25 -1220 45 -1200
rect -175 -1235 45 -1220
rect 80 -1300 100 -1150
rect 310 -1200 380 -1190
rect 310 -1220 325 -1200
rect 365 -1220 380 -1200
rect 310 -1235 380 -1220
rect 5 -1315 40 -1300
rect 5 -1380 10 -1315
rect 35 -1380 40 -1315
rect 5 -1400 40 -1380
rect 65 -1315 100 -1300
rect 65 -1380 70 -1315
rect 95 -1380 100 -1315
rect 65 -1400 100 -1380
rect 255 -1315 290 -1300
rect 255 -1380 260 -1315
rect 285 -1380 290 -1315
rect 255 -1400 290 -1380
rect 315 -1315 350 -1300
rect 315 -1380 320 -1315
rect 345 -1380 350 -1315
rect 315 -1400 350 -1380
rect 255 -1470 275 -1400
rect 85 -1485 275 -1470
rect 85 -1510 105 -1485
rect 215 -1490 275 -1485
rect 215 -1510 230 -1490
rect 85 -1525 230 -1510
rect 410 -1665 450 -1150
rect 525 -1190 610 -200
rect 885 -150 1165 -135
rect 725 -250 795 -240
rect 725 -270 735 -250
rect 775 -270 795 -250
rect 725 -285 795 -270
rect 885 -310 925 -150
rect 1095 -170 1110 -150
rect 1155 -170 1270 -150
rect 1095 -190 1270 -170
rect 1240 -240 1270 -190
rect 1335 -160 1365 -100
rect 1335 -175 1435 -160
rect 1335 -195 1380 -175
rect 1420 -195 1435 -175
rect 1335 -215 1435 -195
rect 1060 -250 1130 -240
rect 1060 -270 1075 -250
rect 1115 -270 1130 -250
rect 1060 -285 1130 -270
rect 1240 -250 1310 -240
rect 1240 -270 1250 -250
rect 1290 -270 1310 -250
rect 1240 -285 1310 -270
rect 885 -330 1095 -310
rect 885 -350 925 -330
rect 1070 -350 1095 -330
rect 1335 -350 1365 -215
rect 755 -365 790 -350
rect 755 -430 760 -365
rect 785 -430 790 -365
rect 755 -450 790 -430
rect 815 -365 925 -350
rect 815 -430 820 -365
rect 845 -375 925 -365
rect 1005 -365 1040 -350
rect 845 -430 850 -375
rect 815 -450 850 -430
rect 1005 -430 1010 -365
rect 1035 -430 1040 -365
rect 1005 -450 1040 -430
rect 1065 -365 1100 -350
rect 1065 -430 1070 -365
rect 1095 -430 1100 -365
rect 1065 -450 1100 -430
rect 1270 -365 1305 -350
rect 1270 -430 1275 -365
rect 1300 -430 1305 -365
rect 1270 -450 1305 -430
rect 1330 -365 1365 -350
rect 1330 -430 1335 -365
rect 1360 -430 1365 -365
rect 1330 -450 1365 -430
rect 760 -525 785 -450
rect 1005 -520 1025 -450
rect 835 -525 1025 -520
rect 760 -535 1025 -525
rect 760 -555 855 -535
rect 835 -560 855 -555
rect 965 -540 1025 -535
rect 1275 -525 1300 -450
rect 1350 -525 1495 -520
rect 1275 -535 1495 -525
rect 965 -560 980 -540
rect 1275 -555 1370 -535
rect 835 -575 980 -560
rect 1350 -560 1370 -555
rect 1480 -560 1495 -535
rect 1350 -575 1495 -560
rect 785 -715 1035 -700
rect 785 -775 820 -715
rect 715 -780 820 -775
rect 1010 -780 1035 -715
rect 1305 -715 1555 -700
rect 1305 -775 1340 -715
rect 715 -800 1035 -780
rect 1235 -780 1340 -775
rect 1530 -780 1555 -715
rect 1235 -800 1555 -780
rect 715 -850 735 -800
rect 1235 -850 1255 -800
rect 695 -865 775 -850
rect 695 -1040 705 -865
rect 765 -1040 775 -865
rect 695 -1050 775 -1040
rect 800 -855 880 -850
rect 945 -855 1025 -850
rect 800 -865 1025 -855
rect 800 -1040 810 -865
rect 870 -905 955 -865
rect 870 -1040 880 -905
rect 800 -1050 880 -1040
rect 945 -1040 955 -905
rect 1015 -1040 1025 -865
rect 945 -1050 1025 -1040
rect 1050 -865 1130 -850
rect 1050 -1040 1060 -865
rect 1120 -1040 1130 -865
rect 1050 -1050 1130 -1040
rect 1215 -865 1295 -850
rect 1215 -1040 1225 -865
rect 1285 -1040 1295 -865
rect 1215 -1050 1295 -1040
rect 1320 -865 1400 -850
rect 1320 -1040 1330 -865
rect 1390 -1040 1400 -865
rect 1320 -1050 1400 -1040
rect 1075 -1070 1115 -1050
rect 870 -1100 1115 -1070
rect 1325 -1100 1355 -1050
rect 525 -1200 780 -1190
rect 525 -1220 720 -1200
rect 760 -1220 780 -1200
rect 525 -1235 780 -1220
rect 870 -1260 910 -1100
rect 1075 -1115 1145 -1100
rect 1325 -1115 1425 -1100
rect 1075 -1135 1090 -1115
rect 1130 -1135 1265 -1115
rect 1075 -1155 1265 -1135
rect 1230 -1190 1265 -1155
rect 1325 -1135 1370 -1115
rect 1410 -1135 1425 -1115
rect 1325 -1155 1425 -1135
rect 1045 -1200 1115 -1190
rect 1045 -1220 1060 -1200
rect 1100 -1220 1115 -1200
rect 1045 -1235 1115 -1220
rect 1230 -1200 1300 -1190
rect 1230 -1220 1240 -1200
rect 1280 -1220 1300 -1200
rect 1230 -1235 1300 -1220
rect 870 -1280 1080 -1260
rect 870 -1300 910 -1280
rect 1055 -1300 1080 -1280
rect 1325 -1300 1355 -1155
rect 740 -1315 775 -1300
rect 740 -1380 745 -1315
rect 770 -1380 775 -1315
rect 740 -1400 775 -1380
rect 800 -1315 910 -1300
rect 800 -1380 805 -1315
rect 830 -1325 910 -1315
rect 990 -1315 1025 -1300
rect 830 -1380 835 -1325
rect 800 -1400 835 -1380
rect 990 -1380 995 -1315
rect 1020 -1380 1025 -1315
rect 990 -1400 1025 -1380
rect 1050 -1315 1085 -1300
rect 1050 -1380 1055 -1315
rect 1080 -1380 1085 -1315
rect 1050 -1400 1085 -1380
rect 1260 -1315 1295 -1300
rect 1260 -1380 1265 -1315
rect 1290 -1380 1295 -1315
rect 1260 -1400 1295 -1380
rect 1320 -1315 1355 -1300
rect 1320 -1380 1325 -1315
rect 1350 -1380 1355 -1315
rect 1320 -1400 1355 -1380
rect 745 -1475 770 -1400
rect 990 -1470 1010 -1400
rect 820 -1475 1010 -1470
rect 745 -1485 1010 -1475
rect 745 -1505 840 -1485
rect 820 -1510 840 -1505
rect 950 -1490 1010 -1485
rect 1265 -1475 1290 -1400
rect 1340 -1475 1485 -1470
rect 1265 -1485 1485 -1475
rect 950 -1510 965 -1490
rect 1265 -1505 1360 -1485
rect 820 -1525 965 -1510
rect 1340 -1510 1360 -1505
rect 1470 -1510 1485 -1485
rect 1340 -1525 1485 -1510
rect 35 -1710 285 -1695
rect 410 -1705 550 -1665
rect 35 -1770 70 -1710
rect -35 -1775 70 -1770
rect 260 -1775 285 -1710
rect -35 -1795 285 -1775
rect -35 -1845 -15 -1795
rect -55 -1860 25 -1845
rect -55 -2035 -45 -1860
rect 15 -2035 25 -1860
rect -55 -2045 25 -2035
rect 50 -1850 130 -1845
rect 195 -1850 275 -1845
rect 50 -1860 275 -1850
rect 50 -2035 60 -1860
rect 120 -1900 205 -1860
rect 120 -2035 130 -1900
rect 50 -2045 130 -2035
rect 195 -2035 205 -1900
rect 265 -2035 275 -1860
rect 195 -2045 275 -2035
rect 300 -1860 380 -1845
rect 300 -2035 310 -1860
rect 370 -2035 380 -1860
rect 300 -2045 380 -2035
rect 325 -2065 365 -2045
rect 120 -2095 365 -2065
rect -40 -2195 30 -2185
rect -40 -2215 -30 -2195
rect 10 -2215 30 -2195
rect -40 -2230 30 -2215
rect 120 -2255 160 -2095
rect 325 -2110 395 -2095
rect 325 -2130 340 -2110
rect 380 -2130 395 -2110
rect 325 -2150 395 -2130
rect 485 -2185 550 -1705
rect 705 -1710 955 -1695
rect 705 -1770 740 -1710
rect 635 -1775 740 -1770
rect 930 -1775 955 -1710
rect 1365 -1710 1615 -1695
rect 1365 -1770 1400 -1710
rect 635 -1795 955 -1775
rect 1295 -1775 1400 -1770
rect 1590 -1775 1615 -1710
rect 1295 -1795 1615 -1775
rect 635 -1845 655 -1795
rect 875 -1845 895 -1795
rect 1295 -1845 1315 -1795
rect 615 -1860 695 -1845
rect 615 -2035 625 -1860
rect 685 -2035 695 -1860
rect 615 -2045 695 -2035
rect 720 -1860 800 -1845
rect 720 -2035 730 -1860
rect 790 -2035 800 -1860
rect 720 -2045 800 -2035
rect 865 -1860 945 -1845
rect 865 -2035 875 -1860
rect 935 -2035 945 -1860
rect 865 -2045 945 -2035
rect 970 -1860 1050 -1845
rect 970 -2035 980 -1860
rect 1040 -2035 1050 -1860
rect 970 -2045 1050 -2035
rect 1275 -1860 1355 -1845
rect 1275 -2035 1285 -1860
rect 1345 -2035 1355 -1860
rect 1275 -2045 1355 -2035
rect 1380 -1860 1460 -1845
rect 1380 -2035 1390 -1860
rect 1450 -2035 1460 -1860
rect 1380 -2045 1460 -2035
rect 735 -2096 780 -2045
rect 981 -2090 1023 -2045
rect 981 -2094 1025 -2090
rect 856 -2096 1025 -2094
rect 735 -2100 1025 -2096
rect 735 -2105 1090 -2100
rect 735 -2125 1035 -2105
rect 1075 -2125 1320 -2105
rect 735 -2145 1320 -2125
rect 295 -2195 365 -2185
rect 295 -2215 310 -2195
rect 350 -2215 365 -2195
rect 295 -2230 365 -2215
rect 485 -2195 700 -2185
rect 485 -2215 640 -2195
rect 680 -2215 700 -2195
rect 485 -2230 700 -2215
rect 120 -2275 330 -2255
rect 120 -2295 160 -2275
rect 305 -2295 330 -2275
rect 735 -2295 755 -2145
rect 1290 -2185 1320 -2145
rect 1385 -2110 1415 -2045
rect 1385 -2125 1485 -2110
rect 1385 -2145 1430 -2125
rect 1470 -2145 1485 -2125
rect 1385 -2165 1485 -2145
rect 965 -2195 1035 -2185
rect 965 -2215 980 -2195
rect 1020 -2215 1035 -2195
rect 965 -2230 1035 -2215
rect 1290 -2195 1360 -2185
rect 1290 -2215 1300 -2195
rect 1340 -2215 1360 -2195
rect 1290 -2230 1360 -2215
rect 1385 -2295 1415 -2165
rect -10 -2310 25 -2295
rect -10 -2375 -5 -2310
rect 20 -2375 25 -2310
rect -10 -2395 25 -2375
rect 50 -2310 160 -2295
rect 50 -2375 55 -2310
rect 80 -2320 160 -2310
rect 240 -2310 275 -2295
rect 80 -2375 85 -2320
rect 50 -2395 85 -2375
rect 240 -2375 245 -2310
rect 270 -2375 275 -2310
rect 240 -2395 275 -2375
rect 300 -2310 335 -2295
rect 300 -2375 305 -2310
rect 330 -2375 335 -2310
rect 300 -2395 335 -2375
rect 660 -2310 695 -2295
rect 660 -2375 665 -2310
rect 690 -2375 695 -2310
rect 660 -2395 695 -2375
rect 720 -2310 755 -2295
rect 720 -2375 725 -2310
rect 750 -2375 755 -2310
rect 720 -2395 755 -2375
rect 910 -2310 945 -2295
rect 910 -2375 915 -2310
rect 940 -2375 945 -2310
rect 910 -2395 945 -2375
rect 970 -2310 1005 -2295
rect 970 -2375 975 -2310
rect 1000 -2375 1005 -2310
rect 970 -2395 1005 -2375
rect 1320 -2310 1355 -2295
rect 1320 -2375 1325 -2310
rect 1350 -2375 1355 -2310
rect 1320 -2395 1355 -2375
rect 1380 -2310 1415 -2295
rect 1380 -2375 1385 -2310
rect 1410 -2375 1415 -2310
rect 1380 -2395 1415 -2375
rect -5 -2470 20 -2395
rect 240 -2465 260 -2395
rect 910 -2465 930 -2395
rect 70 -2470 260 -2465
rect -5 -2480 260 -2470
rect -5 -2500 90 -2480
rect 70 -2505 90 -2500
rect 200 -2485 260 -2480
rect 740 -2480 930 -2465
rect 200 -2505 215 -2485
rect 70 -2520 215 -2505
rect 740 -2505 760 -2480
rect 870 -2485 930 -2480
rect 1325 -2470 1350 -2395
rect 1400 -2470 1545 -2465
rect 1325 -2480 1545 -2470
rect 870 -2505 885 -2485
rect 1325 -2500 1420 -2480
rect 740 -2520 885 -2505
rect 1400 -2505 1420 -2500
rect 1530 -2505 1545 -2480
rect 1400 -2520 1545 -2505
<< viali >>
rect 85 170 275 235
rect 835 170 1025 235
rect 1350 170 1540 235
rect 380 -180 425 -160
rect -15 -270 25 -250
rect 325 -270 365 -250
rect 10 -430 35 -365
rect 320 -430 345 -365
rect 105 -560 215 -535
rect 85 -780 275 -715
rect 380 -1130 420 -1110
rect -15 -1220 25 -1200
rect 325 -1220 365 -1200
rect 10 -1380 35 -1315
rect 320 -1380 345 -1315
rect 105 -1510 215 -1485
rect 735 -270 775 -250
rect 1110 -170 1155 -150
rect 1380 -195 1420 -175
rect 1075 -270 1115 -250
rect 1250 -270 1290 -250
rect 855 -560 965 -535
rect 1370 -560 1480 -535
rect 820 -780 1010 -715
rect 1340 -780 1530 -715
rect 720 -1220 760 -1200
rect 1090 -1135 1130 -1115
rect 1370 -1135 1410 -1115
rect 1060 -1220 1100 -1200
rect 1240 -1220 1280 -1200
rect 840 -1510 950 -1485
rect 1360 -1510 1470 -1485
rect 70 -1775 260 -1710
rect -30 -2215 10 -2195
rect 340 -2130 380 -2110
rect 740 -1775 930 -1710
rect 1400 -1775 1590 -1710
rect 1035 -2125 1075 -2105
rect 310 -2215 350 -2195
rect 640 -2215 680 -2195
rect 1430 -2145 1470 -2125
rect 980 -2215 1020 -2195
rect 1300 -2215 1340 -2195
rect 665 -2375 690 -2310
rect 975 -2375 1000 -2310
rect 90 -2505 200 -2480
rect 760 -2505 870 -2480
rect 1420 -2505 1530 -2480
<< metal1 >>
rect -550 235 1565 250
rect -550 170 85 235
rect 275 170 835 235
rect 1025 170 1350 235
rect 1540 170 1565 235
rect -550 150 1565 170
rect -550 -700 -455 150
rect 365 -160 980 -145
rect 365 -180 380 -160
rect 425 -180 980 -160
rect 365 -200 980 -180
rect 1095 -150 1165 -135
rect 1095 -170 1110 -150
rect 1155 -170 1165 -150
rect 1095 -190 1165 -170
rect 1365 -175 1435 -160
rect 945 -240 980 -200
rect 1365 -195 1380 -175
rect 1420 -195 1435 -175
rect 1365 -215 1435 -195
rect -25 -250 45 -240
rect -25 -270 -15 -250
rect 25 -270 45 -250
rect -25 -285 45 -270
rect 310 -250 380 -240
rect 310 -270 325 -250
rect 365 -270 380 -250
rect 310 -285 380 -270
rect 725 -250 795 -240
rect 725 -270 735 -250
rect 775 -270 795 -250
rect 725 -285 795 -270
rect 945 -250 1130 -240
rect 945 -270 1075 -250
rect 1115 -270 1130 -250
rect 945 -285 1130 -270
rect 1240 -250 1310 -240
rect 1240 -270 1250 -250
rect 1290 -270 1310 -250
rect 1240 -285 1310 -270
rect 5 -365 350 -350
rect 5 -430 10 -365
rect 35 -375 320 -365
rect 35 -430 40 -375
rect 5 -450 40 -430
rect 315 -430 320 -375
rect 345 -430 350 -365
rect 315 -450 350 -430
rect 85 -530 230 -520
rect 85 -560 105 -530
rect 215 -560 230 -530
rect 85 -575 230 -560
rect 835 -530 980 -520
rect 835 -560 855 -530
rect 965 -560 980 -530
rect 835 -575 980 -560
rect 1350 -530 1495 -520
rect 1350 -560 1370 -530
rect 1480 -560 1495 -530
rect 1350 -575 1495 -560
rect -550 -715 1555 -700
rect -550 -780 85 -715
rect 275 -780 820 -715
rect 1010 -780 1340 -715
rect 1530 -780 1555 -715
rect -550 -800 1555 -780
rect -550 -1695 -465 -800
rect 365 -1110 435 -1095
rect 365 -1130 380 -1110
rect 420 -1130 435 -1110
rect 365 -1150 435 -1130
rect 1075 -1115 1145 -1100
rect 1075 -1135 1090 -1115
rect 1130 -1135 1145 -1115
rect 1075 -1155 1145 -1135
rect 1355 -1115 1425 -1100
rect 1355 -1135 1370 -1115
rect 1410 -1135 1425 -1115
rect 1355 -1155 1425 -1135
rect -25 -1200 45 -1190
rect -25 -1220 -15 -1200
rect 25 -1220 45 -1200
rect -25 -1235 45 -1220
rect 310 -1200 380 -1190
rect 310 -1220 325 -1200
rect 365 -1220 380 -1200
rect 310 -1235 380 -1220
rect 710 -1200 780 -1190
rect 710 -1220 720 -1200
rect 760 -1220 780 -1200
rect 710 -1235 780 -1220
rect 1045 -1200 1115 -1190
rect 1045 -1220 1060 -1200
rect 1100 -1220 1115 -1200
rect 1045 -1235 1115 -1220
rect 1230 -1200 1300 -1190
rect 1230 -1220 1240 -1200
rect 1280 -1220 1300 -1200
rect 1230 -1235 1300 -1220
rect 5 -1315 350 -1300
rect 5 -1380 10 -1315
rect 35 -1325 320 -1315
rect 35 -1380 40 -1325
rect 5 -1400 40 -1380
rect 315 -1380 320 -1325
rect 345 -1380 350 -1315
rect 315 -1400 350 -1380
rect 85 -1480 230 -1470
rect 85 -1510 105 -1480
rect 215 -1510 230 -1480
rect 85 -1525 230 -1510
rect 820 -1480 965 -1470
rect 820 -1510 840 -1480
rect 950 -1510 965 -1480
rect 820 -1525 965 -1510
rect 1340 -1480 1485 -1470
rect 1340 -1510 1360 -1480
rect 1470 -1510 1485 -1480
rect 1340 -1525 1485 -1510
rect -550 -1710 1615 -1695
rect -550 -1775 70 -1710
rect 260 -1775 740 -1710
rect 930 -1775 1400 -1710
rect 1590 -1775 1615 -1710
rect -550 -1795 1615 -1775
rect -550 -1800 -95 -1795
rect 325 -2100 395 -2095
rect 325 -2110 870 -2100
rect 325 -2130 340 -2110
rect 380 -2130 870 -2110
rect 325 -2150 870 -2130
rect 1020 -2105 1090 -2100
rect 1020 -2125 1035 -2105
rect 1075 -2125 1090 -2105
rect 1020 -2145 1090 -2125
rect 1415 -2125 1485 -2110
rect 1415 -2145 1430 -2125
rect 1470 -2145 1485 -2125
rect 830 -2185 870 -2150
rect 1415 -2165 1485 -2145
rect -40 -2195 30 -2185
rect -40 -2215 -30 -2195
rect 10 -2215 30 -2195
rect -40 -2230 30 -2215
rect 295 -2195 365 -2185
rect 295 -2215 310 -2195
rect 350 -2215 365 -2195
rect 295 -2230 365 -2215
rect 630 -2195 700 -2185
rect 630 -2215 640 -2195
rect 680 -2215 700 -2195
rect 630 -2230 700 -2215
rect 830 -2195 1035 -2185
rect 830 -2215 980 -2195
rect 1020 -2215 1035 -2195
rect 830 -2230 1035 -2215
rect 1290 -2195 1360 -2185
rect 1290 -2215 1300 -2195
rect 1340 -2215 1360 -2195
rect 1290 -2230 1360 -2215
rect 660 -2310 1005 -2295
rect 660 -2375 665 -2310
rect 690 -2320 975 -2310
rect 690 -2375 695 -2320
rect 660 -2395 695 -2375
rect 970 -2375 975 -2320
rect 1000 -2375 1005 -2310
rect 970 -2395 1005 -2375
rect 70 -2475 215 -2465
rect 70 -2505 90 -2475
rect 200 -2505 215 -2475
rect 70 -2520 215 -2505
rect 740 -2475 885 -2465
rect 740 -2505 760 -2475
rect 870 -2505 885 -2475
rect 740 -2520 885 -2505
rect 1400 -2475 1545 -2465
rect 1400 -2505 1420 -2475
rect 1530 -2505 1545 -2475
rect 1400 -2520 1545 -2505
<< via1 >>
rect 105 -535 215 -530
rect 105 -560 215 -535
rect 855 -535 965 -530
rect 855 -560 965 -535
rect 1370 -535 1480 -530
rect 1370 -560 1480 -535
rect 105 -1485 215 -1480
rect 105 -1510 215 -1485
rect 840 -1485 950 -1480
rect 840 -1510 950 -1485
rect 1360 -1485 1470 -1480
rect 1360 -1510 1470 -1485
rect 90 -2480 200 -2475
rect 90 -2505 200 -2480
rect 760 -2480 870 -2475
rect 760 -2505 870 -2480
rect 1420 -2480 1530 -2475
rect 1420 -2505 1530 -2480
<< metal2 >>
rect -370 -530 1495 -520
rect -370 -560 105 -530
rect 215 -560 855 -530
rect 965 -560 1370 -530
rect 1480 -560 1495 -530
rect -370 -575 1495 -560
rect -370 -1470 -300 -575
rect -370 -1480 1485 -1470
rect -370 -1510 105 -1480
rect 215 -1510 840 -1480
rect 950 -1510 1360 -1480
rect 1470 -1510 1485 -1480
rect -370 -1525 1485 -1510
rect -370 -2465 -300 -1525
rect -370 -2475 1545 -2465
rect -370 -2505 90 -2475
rect 200 -2505 760 -2475
rect 870 -2505 1420 -2475
rect 1530 -2505 1545 -2475
rect -370 -2520 1545 -2505
<< labels >>
rlabel metal1 -200 200 -200 200 1 vdd
port 1 n
rlabel metal2 -145 -2485 -145 -2485 1 gnd
port 2 n
rlabel metal1 -15 -280 -15 -280 1 l(i-1)
port 3 n
rlabel metal1 355 -280 355 -280 1 l(x-1)
port 4 n
rlabel metal1 365 -1230 365 -1230 1 cl(i-2)
port 5 n
rlabel metal1 -15 -2225 -15 -2225 1 l(y-1)
port 6 n
rlabel metal1 355 -2220 355 -2220 1 l(z-1)
port 7 n
rlabel metal1 785 -275 785 -275 1 l(i)
port 8 n
rlabel metal1 1105 -1230 1105 -1230 1 cl(i-1)
port 9 n
rlabel metal1 1095 -1150 1095 -1150 1 l(y)
port 11 n
rlabel metal1 1125 -180 1125 -180 1 l(x)
port 12 n
rlabel metal1 1405 -205 1405 -205 1 l(x)
port 13 n
rlabel metal1 1400 -1150 1400 -1150 1 l(y)
port 14 n
rlabel metal1 1440 -2160 1440 -2160 1 l(z)
port 15 n
rlabel metal1 1045 -2140 1045 -2140 1 l(z)
port 15 n
<< end >>
